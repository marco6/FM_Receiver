--test bench loop filter
--mohamed ali version