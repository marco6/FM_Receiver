--test bench loop filter
