--test bench loop filter

entity test_loopFilter is
end entity;

architecture Behavioral of test_loopFilter is
begin
 -- TODO: this is just to make ghdl happy
end architecture;
