--here the code of loop filter
--